//***********************************************
//Project Name               :
//File Name                  :
//Author                     :ZJL
//Date of Creation           :20190920
//Functional Description     :图像数据仿真
//
//Revision History           :
//Change Log                 :
//***********************************************
`timescale 1ns / 1ns
// `include "../../rtl/ghe_include.v"
module tb;
        // auto generated by tools/config_tb.py
        parameter PIXEL_CLK = 40;  //100MHz
        parameter CLK_PERIOD = 1000 / PIXEL_CLK;  //像素时钟周期-10ns
        parameter FRAME_RATE = 50;  //帧频
        parameter WIDTH =10'd640;  //分辨率：宽度
        parameter LINE_BLANK = 100;  //行消隐期
        parameter TOTAL_COL = (WIDTH + LINE_BLANK);  //每行总像素数-740
        parameter HIDTH = 10'd512;  //分辨率：高度
        parameter EXTRA_LINES = 0;  //多输出的行数
        parameter TOTAL_ROW = (HIDTH + EXTRA_LINES);  //总行数-1034
        parameter TOTAL_PIXEL = TOTAL_COL * TOTAL_ROW;  //每帧总像素数
        parameter FRAME_PERIOD = 1_000_000_000 / FRAME_RATE;  //帧周期-16,666,666.66666667ns
        parameter VIDEO_BEGIN = 100;//(PIXEL_CLK * 1_000_000 / FRAME_RATE - (TOTAL_COL * TOTAL_ROW)) / 2;  //1帧内总时钟数-总像素数
        parameter CNT_FIELD = PIXEL_CLK * 1_000_000 / FRAME_RATE;  //帧同步计数
        parameter DW = 16;  //数据宽度
        parameter CW = 10;  //地址宽度
        // generated end                                                                                                                                                                                                                                                                                                                                                                                                                                            
    parameter IMAGE_WIDTH = WIDTH;
    parameter IMAGE_HEIGHT = HIDTH;
    //信号列表
    reg                  rst_n;  //reset @high voltage

    wire                 i_clk;  //clock
    wire                 i_rst_n;  //reset @high voltage
    wire                 i_clk_mul4;  //clock
    reg                  sys_clk_x4;  //reset @high voltage
    wire                 i_mul4_rst_n;  //reset @high voltage

    reg                  in_pulse;  //input signal
    wire    [       7:0] o_data;  //data after scale
    wire                 o_dvalid;  //data valid after scale
    reg     [    DW-1:0] data_tmp;
    wire    [     1-1:0] data_tmp2_vld;
    reg     [    DW-1:0] data_tmp2;
    wire    [     1-1:0] h_valid_dly;
    wire    [    DW-1:0] data_tmp_dly;
    integer              addr;  //memory address

    reg     [     1-1:0] field_sync;
    wire    [     1-1:0] field_rst;
    reg     [    32-1:0] cnt_field_sync;
    wire    [     1-1:0] wait_time_add;
    reg     [     1-1:0] en_cnt_wait_time;
    reg     [    32-1:0] cnt_wait_time;
    wire    [     1-1:0] wait_done;
    reg     [     1-1:0] flag_image;
    reg     [    12-1:0] hcnt;
    reg     [    12-1:0] vcnt;
    wire    [     1-1:0] h_valid;
    wire    [     1-1:0] v_valid;

    wire                 i_Sys_clk;
    wire                 i_Rst_n;
    wire                 aresetn;
    wire    [1  - 1 : 0] field_rst_neg_delay;
    gen_field_rst #(
        .FIELD_RST_DELAY(200)
    ) u_gen_rst (
        .i_Sys_clk   (i_Sys_clk),
        .i_Rst_n     (i_Rst_n),
        .i_Field_sync(h_valid),
        .o_Field_rst (field_rst_neg_delay)
    );
    //**********************************************************************************************
    //系统时钟   
    // initial begin
    //     sys_clk = 0;
    //     forever #(CLK_PERIOD / 2) sys_clk = ~sys_clk;
    // end

    // parameter PIXEL_CLK = 10;  //50MHz
    parameter PIXEL_CLK_x4 = PIXEL_CLK * 4;  //50MHz
    parameter CLKx4_PERIOD = 1000 / PIXEL_CLK_x4;  //像素时钟周期-20ns
    reg  [1:0] clk_div;
    wire       sys_clk;
    initial begin
        sys_clk_x4 = 0;
        forever #(CLKx4_PERIOD / 2) sys_clk_x4 = ~sys_clk_x4;
    end
    always @(posedge sys_clk_x4) begin
        if (~i_Rst_n) begin
            clk_div <= 2'b00;
        end else if (clk_div == 2'b11) begin
            clk_div <= 2'b00;
        end else begin
            clk_div <= clk_div + 1'b1;
        end
    end

    assign sys_clk      = (clk_div == 2'b11 || clk_div < 2'b01) ? 1'b1 : 1'b0;


    assign aresetn      = rst_n;
    assign i_Sys_clk    = sys_clk;  //sys_clk;
    assign i_Rst_n      = rst_n;
    assign i_clk        = sys_clk;  //sys_clk;
    assign i_rst_n      = rst_n;
    assign i_clk_mul4   = sys_clk_x4;
    assign i_mul4_rst_n = rst_n;
    wire axi_aclk      ;assign axi_aclk     =  i_clk_mul4   ;
    wire axi_aresetn   ;assign axi_aresetn  =  i_mul4_rst_n ;
    //*********************************************行场同步信号*************************************************
    // 帧同步信号产生
    always @(posedge i_Sys_clk) begin
        if (~i_Rst_n) begin
            cnt_field_sync <= 'd0;
        end else if (cnt_field_sync == CNT_FIELD - 1) begin
            cnt_field_sync <= 'd0;
        end else begin
            cnt_field_sync <= cnt_field_sync + 'd1;
        end
    end
    always @(posedge i_Sys_clk) begin
        if (~i_Rst_n) begin
            field_sync <= 'd1;
        end else if (cnt_field_sync == CNT_FIELD - 1) begin
            field_sync <= ~field_sync;
        end else begin
            field_sync <= field_sync;
        end
    end
    assign field_rst     = cnt_field_sync == 1;  //CNT_FIELD-1
    //------------------行计数-----------------------
    assign wait_time_add = field_rst;
    always @(posedge sys_clk) begin
        if (~rst_n) begin
            cnt_wait_time <= 'd0;
        end else if (en_cnt_wait_time) begin  //只有在有效才计数
            cnt_wait_time <= cnt_wait_time + 'd1;
        end else begin
            cnt_wait_time <= 'd0;
        end
    end

    always @(posedge sys_clk) begin
        if (~rst_n) begin
            en_cnt_wait_time <= 'd0;
        end else if (cnt_wait_time == VIDEO_BEGIN - 1) begin  //结束计数条件
            en_cnt_wait_time <= 'd0;
        end else if (field_rst) begin  //开始计数条件
            en_cnt_wait_time <= 'd1;
        end else begin
            en_cnt_wait_time <= en_cnt_wait_time;
        end
    end
    assign wait_done = (cnt_wait_time == VIDEO_BEGIN - 1);

    always @(posedge sys_clk) begin
        if (~rst_n) begin
            flag_image <= 'd0;
        end else if (vcnt == TOTAL_ROW - 1 && hcnt == WIDTH - 1) begin  //结束计数条件
            flag_image <= 'd0;
        end else if (wait_done) begin  //开始计数条件
            flag_image <= 'd1;
        end else begin
            flag_image <= flag_image;
        end
    end
    always @(posedge sys_clk) begin
        if (~rst_n) begin
            hcnt <= 'd0;
        end else if (field_rst_neg_delay) begin
            hcnt <= 0;
        end else if (flag_image) begin  //结束计数条件
            if (hcnt == TOTAL_COL - 1) hcnt <= 'd0;
            else hcnt <= hcnt + 'd1;
        end else begin
            hcnt <= 'd0;
        end
    end
    assign h_valid = (flag_image && hcnt < WIDTH);
    assign v_valid = (flag_image && vcnt < HIDTH);
    always @(posedge sys_clk) begin
        if (~rst_n) begin
            vcnt <= 'd0;
        end else if (field_rst_neg_delay) begin
            vcnt <= 0;
        end else if (flag_image) begin  //结束计数条件
            if (hcnt == TOTAL_COL - 1) vcnt <= vcnt + 'd1;
            else vcnt <= vcnt;
        end else begin
            vcnt <= 'd0;
        end
    end
    //**********************************************************************************************
    //------------------任务------------------------
    //*任务：系统初始化
    task task_sysinit;
        begin
            in_pulse = 0;
        end
    endtask

    //*任务：Generate global reset
    task task_reset;
        begin
            rst_n = 0;
            repeat (2) @(negedge sys_clk_x4);
            rst_n = 1;
        end
    endtask


    //*任务：读取文件到内存
    reg [DW-1:0] reg_mem    [0:WIDTH*HIDTH-1];  //! memory
    reg [DW-1:0] reg_mem0[0:WIDTH*HIDTH-1];
    reg [DW-1:0] reg_mem1[0:WIDTH*HIDTH-1];
    reg [DW-1:0] reg_mem2[0:WIDTH*HIDTH-1];
    reg [DW-1:0] reg_mem3[0:WIDTH*HIDTH-1];
    reg [DW-1:0] reg_mem4[0:WIDTH*HIDTH-1];
    reg [DW-1:0] reg_mem5[0:WIDTH*HIDTH-1];
    reg [DW-1:0] reg_mem6[0:WIDTH*HIDTH-1];
    reg [DW-1:0] reg_mem7[0:WIDTH*HIDTH-1];
    reg [DW-1:0] reg_mem8[0:WIDTH*HIDTH-1];
    reg [DW-1:0] reg_mem9[0:WIDTH*HIDTH-1];
    reg [DW-1:0] reg_mem10[0:WIDTH*HIDTH-1];
    reg [8 -1:0] reg_mem_low[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem11[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem12[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem13[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem14[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem15[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem16[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem17[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem18[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem19[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem20[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem21[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem22[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem23[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem24[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem25[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem26[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem27[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem28[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem29[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem30[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem31[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem32[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem33[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem34[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem35[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem36[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem37[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem38[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem39[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem40[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem41[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem42[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem43[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem44[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem45[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem46[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem47[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem48[0:WIDTH*HIDTH-1];
    // reg [DW-1:0] reg_mem49[0:WIDTH*HIDTH-1];
    task load_data2mem;
        begin
            $readmemh("../output/ghe_in.txt", reg_mem0);
            $readmemh("../output/ghe_in.txt", reg_mem1);
            $readmemh("../output/ghe_in.txt", reg_mem2);
            $readmemh("../output/ghe_in.txt", reg_mem3);
            $readmemh("../output/ghe_in.txt", reg_mem4);
            $readmemh("../output/ghe_in.txt", reg_mem5);
            $readmemh("../output/ghe_in.txt", reg_mem6);
            $readmemh("../output/ghe_in.txt", reg_mem7);
            $readmemh("../output/ghe_in.txt", reg_mem8);
            $readmemh("../output/ghe_in.txt", reg_mem9);
            $readmemh("../output/ghe_in.txt", reg_mem10);
            $readmemh("../output/ghe_out.txt", reg_mem_low);
        end
    endtask

    //-----------------存储器地址------------------------
    reg [8  - 1 : 0] frame_num;
    always @(posedge i_Sys_clk) begin
        if (~i_Rst_n) begin
            frame_num <= 'd0;
        end else if (field_rst) begin
            frame_num <= frame_num + 'd1;
        end else begin
            frame_num <= frame_num;
        end
    end
    
    always @(posedge i_Sys_clk) begin
        if (field_rst) begin
            $display("******************* frame_num = %d", frame_num);
        end
    end
    //生成存储器地址
    always @(posedge sys_clk) begin
        if (!rst_n) begin
            addr <= 0;
        end else if (field_rst_neg_delay) begin
            addr <= 0;
        end else if (h_valid) begin
            addr <= addr + 1;
        end
    end
    
    always @(*) begin
        if (!rst_n) begin
            data_tmp <= 0;
            data_tmp2 <= 0;
        end else begin
            case (frame_num - 'd1)
                0: begin
                    data_tmp     <= reg_mem0[addr];
                    data_tmp2     <= reg_mem_low[addr];
                end  //reg_mem0[addr];
                1: begin
                    data_tmp     <= reg_mem1[addr];
                    data_tmp2     <= reg_mem_low[addr];
                end  //reg_mem1[addr];
                2: begin
                    data_tmp     <= reg_mem2[addr];
                    data_tmp2     <= reg_mem_low[addr];
                end  //reg_mem2[addr];
                3: begin
                    data_tmp     <= reg_mem3[addr];
                    data_tmp2     <= reg_mem_low[addr];
                end  //reg_mem2[addr];
                4: begin
                    data_tmp     <= reg_mem4[addr];
                    data_tmp2     <= reg_mem_low[addr];
                end  //reg_mem2[addr];
                5: begin
                    data_tmp     <= reg_mem5[addr];
                    data_tmp2     <= reg_mem_low[addr];
                end  //reg_mem2[addr];
                6: begin
                    data_tmp     <= reg_mem6[addr];
                    data_tmp2     <= reg_mem_low[addr];
                end  //reg_mem2[addr];
                7: begin
                    data_tmp     <= reg_mem7[addr];
                    data_tmp2     <= reg_mem_low[addr];
                end  //reg_mem2[addr];
                8: begin
                    data_tmp     <= reg_mem8[addr];
                    data_tmp2     <= reg_mem_low[addr];
                end  //reg_mem2[addr];
                9: begin
                    data_tmp     <= reg_mem9[addr];
                    data_tmp2     <= reg_mem_low[addr];
                end  //reg_mem2[addr];
                10: begin
                    data_tmp     <= reg_mem10[addr];
                    data_tmp2     <= reg_mem_low[addr];
                end  //reg_mem2[addr];
                default: ;
            endcase
        end
    end
    //----------------------系统初始化------------------------
    initial begin
        task_sysinit;
        task_reset;
        load_data2mem;

        #100 @(posedge sys_clk) in_pulse = 1;
        @(posedge sys_clk) in_pulse = 0;
        // #10000000;
        // #20;
        // $stop;
    end
    assign data_tmp2_vld = h_valid;
    //**********************************************************************************************

    `define S0_NUMBER 0
    `define S1_NUMBER 1
    `define M0_NUMBER 2
    localparam                          DVP_DATA_WIDTH            = 16   ;
    localparam                          AXI_DW                    = 32;//256   ;
    localparam                          AXI_AW                    = 32    ;
    localparam                          AXI_ID_WIDTH              = 8     ;
    localparam                          AXI_SW                    = AXI_DW / 8;

    localparam S_COUNT = 2;
    localparam M_COUNT = 1;
    localparam AXI_CNT = S_COUNT + M_COUNT;

    wire               [1              - 1 : 0]user0_wr_rst      ;
    wire               [1              - 1 : 0]user0_wr_clk      ;
    wire               [1              - 1 : 0]user0_wr_vs       ;
    wire               [1              - 1 : 0]user0_wr_hs       ;
    wire               [DVP_DATA_WIDTH - 1 : 0]user0_wr_data     ;
    wire               [AXI_AW         - 1 : 0]user0_wr_axi_addr ;
    wire               [1              - 1 : 0]user1_wr_rst      ;
    wire               [1              - 1 : 0]user1_wr_clk      ;
    wire               [1              - 1 : 0]user1_wr_vs       ;
    wire               [1              - 1 : 0]user1_wr_hs       ;
    wire               [DVP_DATA_WIDTH - 1 : 0]user1_wr_data     ;
    wire               [AXI_AW         - 1 : 0]user1_wr_axi_addr ;
    wire               [1              - 1 : 0]user0_rd_rst      ;
    wire               [1              - 1 : 0]user0_rd_clk      ;
    wire               [1              - 1 : 0]user0_rd_vs       ;
    wire               [1              - 1 : 0]user0_rd_hs       ;
    wire               [DVP_DATA_WIDTH - 1 : 0]user0_rd_data     ;
    wire               [AXI_AW         - 1 : 0]user0_rd_axi_addr ;
    wire               [1              - 1 : 0]user1_rd_rst      ;
    wire               [1              - 1 : 0]user1_rd_clk      ;
    wire               [1              - 1 : 0]user1_rd_vs       ;
    wire               [1              - 1 : 0]user1_rd_hs       ;
    wire               [DVP_DATA_WIDTH - 1 : 0]user1_rd_data     ;
    wire               [AXI_AW         - 1 : 0]user1_rd_axi_addr ;

    assign user0_wr_clk =  i_clk        ;
    assign user1_wr_clk =  i_clk        ;
    assign user0_rd_clk =  i_clk        ;
    assign user1_rd_clk =  i_clk        ;
    // assign user0_wr_rst =  field_rst_neg_delay        ;
    // assign user0_rd_rst =  field_rst_neg_delay        ;
    // assign user1_wr_rst =  field_rst_neg_delay        ;
    // assign user1_rd_rst =  field_rst_neg_delay        ;
    wire [          AXI_CNT*8-1:0] axi_awid;
    wire [     AXI_CNT*AXI_AW-1:0] axi_awaddr;
    wire [          AXI_CNT*8-1:0] axi_awlen;
    wire [          AXI_CNT*3-1:0] axi_awsize;
    wire [          AXI_CNT*2-1:0] axi_awburst;
    wire [            AXI_CNT-1:0] axi_awlock;
    wire [          AXI_CNT*4-1:0] axi_awcache;
    wire [          AXI_CNT*3-1:0] axi_awprot;
    wire [            AXI_CNT-1:0] axi_awvalid;
    wire [            AXI_CNT-1:0] axi_awready;
    wire [     AXI_CNT*AXI_DW-1:0] axi_wdata;
    wire [     AXI_CNT*AXI_SW-1:0] axi_wstrb;
    wire [            AXI_CNT-1:0] axi_wlast;
    wire [            AXI_CNT-1:0] axi_wvalid;
    wire [            AXI_CNT-1:0] axi_wready;
    wire [          AXI_CNT*8-1:0] axi_bid;
    wire [          AXI_CNT*2-1:0] axi_bresp;
    wire [            AXI_CNT-1:0] axi_bvalid;
    wire [            AXI_CNT-1:0] axi_bready;
    wire [          AXI_CNT*8-1:0] axi_arid;
    wire [     AXI_CNT*AXI_AW-1:0] axi_araddr;
    wire [          AXI_CNT*8-1:0] axi_arlen;
    wire [          AXI_CNT*3-1:0] axi_arsize;
    wire [          AXI_CNT*2-1:0] axi_arburst;
    wire [            AXI_CNT-1:0] axi_arlock;
    wire [          AXI_CNT*4-1:0] axi_arcache;
    wire [          AXI_CNT*3-1:0] axi_arprot;
    wire [            AXI_CNT-1:0] axi_arvalid;
    wire [            AXI_CNT-1:0] axi_arready;
    wire [          AXI_CNT*8-1:0] axi_rid;
    wire [     AXI_CNT*AXI_DW-1:0] axi_rdata;
    wire [          AXI_CNT*2-1:0] axi_rresp;
    wire [            AXI_CNT-1:0] axi_rlast;
    wire [            AXI_CNT-1:0] axi_rvalid;
    wire [            AXI_CNT-1:0] axi_rready;
    wire [ 1*8-1      : 0 ] m0_axi_awid     ,s0_axi_awid     ,s1_axi_awid     ;
    wire [ 1*AXI_AW-1 : 0 ] m0_axi_awaddr   ,s0_axi_awaddr   ,s1_axi_awaddr   ;
    wire [ 1*8-1      : 0 ] m0_axi_awlen    ,s0_axi_awlen    ,s1_axi_awlen    ;
    wire [ 1*3-1      : 0 ] m0_axi_awsize   ,s0_axi_awsize   ,s1_axi_awsize   ;
    wire [ 1*2-1      : 0 ] m0_axi_awburst  ,s0_axi_awburst  ,s1_axi_awburst  ;
    wire [ 1-1        : 0 ] m0_axi_awlock   ,s0_axi_awlock   ,s1_axi_awlock   ;
    wire [ 1*4-1      : 0 ] m0_axi_awcache  ,s0_axi_awcache  ,s1_axi_awcache  ;
    wire [ 1*3-1      : 0 ] m0_axi_awprot   ,s0_axi_awprot   ,s1_axi_awprot   ;
    wire [ 1-1        : 0 ] m0_axi_awvalid  ,s0_axi_awvalid  ,s1_axi_awvalid  ;
    wire [ 1-1        : 0 ] m0_axi_awready  ,s0_axi_awready  ,s1_axi_awready  ;
    wire [ 1*AXI_DW-1 : 0 ] m0_axi_wdata    ,s0_axi_wdata    ,s1_axi_wdata    ;
    wire [ 1*AXI_SW-1 : 0 ] m0_axi_wstrb    ,s0_axi_wstrb    ,s1_axi_wstrb    ;
    wire [ 1-1        : 0 ] m0_axi_wlast    ,s0_axi_wlast    ,s1_axi_wlast    ;
    wire [ 1-1        : 0 ] m0_axi_wvalid   ,s0_axi_wvalid   ,s1_axi_wvalid   ;
    wire [ 1-1        : 0 ] m0_axi_wready   ,s0_axi_wready   ,s1_axi_wready   ;
    wire [ 1*8-1      : 0 ] m0_axi_bid      ,s0_axi_bid      ,s1_axi_bid      ;
    wire [ 1*2-1      : 0 ] m0_axi_bresp    ,s0_axi_bresp    ,s1_axi_bresp    ;
    wire [ 1-1        : 0 ] m0_axi_bvalid   ,s0_axi_bvalid   ,s1_axi_bvalid   ;
    wire [ 1-1        : 0 ] m0_axi_bready   ,s0_axi_bready   ,s1_axi_bready   ;
    wire [ 1*8-1      : 0 ] m0_axi_arid     ,s0_axi_arid     ,s1_axi_arid     ;
    wire [ 1*AXI_AW-1 : 0 ] m0_axi_araddr   ,s0_axi_araddr   ,s1_axi_araddr   ;
    wire [ 1*8-1      : 0 ] m0_axi_arlen    ,s0_axi_arlen    ,s1_axi_arlen    ;
    wire [ 1*3-1      : 0 ] m0_axi_arsize   ,s0_axi_arsize   ,s1_axi_arsize   ;
    wire [ 1*2-1      : 0 ] m0_axi_arburst  ,s0_axi_arburst  ,s1_axi_arburst  ;
    wire [ 1-1        : 0 ] m0_axi_arlock   ,s0_axi_arlock   ,s1_axi_arlock   ;
    wire [ 1*4-1      : 0 ] m0_axi_arcache  ,s0_axi_arcache  ,s1_axi_arcache  ;
    wire [ 1*3-1      : 0 ] m0_axi_arprot   ,s0_axi_arprot   ,s1_axi_arprot   ;
    wire [ 1-1        : 0 ] m0_axi_arvalid  ,s0_axi_arvalid  ,s1_axi_arvalid  ;
    wire [ 1-1        : 0 ] m0_axi_arready  ,s0_axi_arready  ,s1_axi_arready  ;
    wire [ 1*8-1      : 0 ] m0_axi_rid      ,s0_axi_rid      ,s1_axi_rid      ;
    wire [ 1*AXI_DW-1 : 0 ] m0_axi_rdata    ,s0_axi_rdata    ,s1_axi_rdata    ;
    wire [ 1*2-1      : 0 ] m0_axi_rresp    ,s0_axi_rresp    ,s1_axi_rresp    ;
    wire [ 1-1        : 0 ] m0_axi_rlast    ,s0_axi_rlast    ,s1_axi_rlast    ;
    wire [ 1-1        : 0 ] m0_axi_rvalid   ,s0_axi_rvalid   ,s1_axi_rvalid   ;
    wire [ 1-1        : 0 ] m0_axi_rready   ,s0_axi_rready   ,s1_axi_rready   ;

    assign m0_axi_awid     = axi_awid    [`M0_NUMBER*8         +: 1*8      ];
    assign m0_axi_awaddr   = axi_awaddr  [`M0_NUMBER*AXI_AW    +: 1*AXI_AW ];
    assign m0_axi_awlen    = axi_awlen   [`M0_NUMBER*8         +: 1*8      ];
    assign m0_axi_awsize   = axi_awsize  [`M0_NUMBER*3         +: 1*3      ];
    assign m0_axi_awburst  = axi_awburst [`M0_NUMBER*2         +: 1*2      ];
    assign m0_axi_awlock   = axi_awlock  [`M0_NUMBER           +: 1        ];
    assign m0_axi_awcache  = axi_awcache [`M0_NUMBER*4         +: 1*4      ];
    assign m0_axi_awprot   = axi_awprot  [`M0_NUMBER*3         +: 1*3      ];
    assign m0_axi_awvalid  = axi_awvalid [`M0_NUMBER           +: 1        ];
    assign m0_axi_awready  = axi_awready [`M0_NUMBER           +: 1        ];
    assign m0_axi_wdata    = axi_wdata   [`M0_NUMBER*AXI_DW    +: 1*AXI_DW ];
    assign m0_axi_wstrb    = axi_wstrb   [`M0_NUMBER*AXI_SW    +: 1*AXI_SW ];
    assign m0_axi_wlast    = axi_wlast   [`M0_NUMBER           +: 1        ];
    assign m0_axi_wvalid   = axi_wvalid  [`M0_NUMBER           +: 1        ];
    assign m0_axi_wready   = axi_wready  [`M0_NUMBER           +: 1        ];
    assign m0_axi_bid      = axi_bid     [`M0_NUMBER*8         +: 1*8      ];
    assign m0_axi_bresp    = axi_bresp   [`M0_NUMBER*2         +: 1*2      ];
    assign m0_axi_bvalid   = axi_bvalid  [`M0_NUMBER           +: 1        ];
    assign m0_axi_bready   = axi_bready  [`M0_NUMBER           +: 1        ];
    assign m0_axi_arid     = axi_arid    [`M0_NUMBER*8         +: 1*8      ];
    assign m0_axi_araddr   = axi_araddr  [`M0_NUMBER*AXI_AW    +: 1*AXI_AW ];
    assign m0_axi_arlen    = axi_arlen   [`M0_NUMBER*8         +: 1*8      ];
    assign m0_axi_arsize   = axi_arsize  [`M0_NUMBER*3         +: 1*3      ];
    assign m0_axi_arburst  = axi_arburst [`M0_NUMBER*2         +: 1*2      ];
    assign m0_axi_arlock   = axi_arlock  [`M0_NUMBER           +: 1        ];
    assign m0_axi_arcache  = axi_arcache [`M0_NUMBER*4         +: 1*4      ];
    assign m0_axi_arprot   = axi_arprot  [`M0_NUMBER*3         +: 1*3      ];
    assign m0_axi_arvalid  = axi_arvalid [`M0_NUMBER           +: 1        ];
    assign m0_axi_arready  = axi_arready [`M0_NUMBER           +: 1        ];
    assign m0_axi_rid      = axi_rid     [`M0_NUMBER*8         +: 1*8      ];
    assign m0_axi_rdata    = axi_rdata   [`M0_NUMBER*AXI_DW    +: 1*AXI_DW ];
    assign m0_axi_rresp    = axi_rresp   [`M0_NUMBER*2         +: 1*2      ];
    assign m0_axi_rlast    = axi_rlast   [`M0_NUMBER           +: 1        ];
    assign m0_axi_rvalid   = axi_rvalid  [`M0_NUMBER           +: 1        ];
    assign m0_axi_rready   = axi_rready  [`M0_NUMBER           +: 1        ];
    assign s0_axi_awid     = axi_awid    [`S0_NUMBER*8         +: 1*8      ];
    assign s0_axi_awaddr   = axi_awaddr  [`S0_NUMBER*AXI_AW    +: 1*AXI_AW ];
    assign s0_axi_awlen    = axi_awlen   [`S0_NUMBER*8         +: 1*8      ];
    assign s0_axi_awsize   = axi_awsize  [`S0_NUMBER*3         +: 1*3      ];
    assign s0_axi_awburst  = axi_awburst [`S0_NUMBER*2         +: 1*2      ];
    assign s0_axi_awlock   = axi_awlock  [`S0_NUMBER           +: 1        ];
    assign s0_axi_awcache  = axi_awcache [`S0_NUMBER*4         +: 1*4      ];
    assign s0_axi_awprot   = axi_awprot  [`S0_NUMBER*3         +: 1*3      ];
    assign s0_axi_awvalid  = axi_awvalid [`S0_NUMBER           +: 1        ];
    assign s0_axi_awready  = axi_awready [`S0_NUMBER           +: 1        ];
    assign s0_axi_wdata    = axi_wdata   [`S0_NUMBER*AXI_DW    +: 1*AXI_DW ];
    assign s0_axi_wstrb    = axi_wstrb   [`S0_NUMBER*AXI_SW    +: 1*AXI_SW ];
    assign s0_axi_wlast    = axi_wlast   [`S0_NUMBER           +: 1        ];
    assign s0_axi_wvalid   = axi_wvalid  [`S0_NUMBER           +: 1        ];
    assign s0_axi_wready   = axi_wready  [`S0_NUMBER           +: 1        ];
    assign s0_axi_bid      = axi_bid     [`S0_NUMBER*8         +: 1*8      ];
    assign s0_axi_bresp    = axi_bresp   [`S0_NUMBER*2         +: 1*2      ];
    assign s0_axi_bvalid   = axi_bvalid  [`S0_NUMBER           +: 1        ];
    assign s0_axi_bready   = axi_bready  [`S0_NUMBER           +: 1        ];
    assign s0_axi_arid     = axi_arid    [`S0_NUMBER*8         +: 1*8      ];
    assign s0_axi_araddr   = axi_araddr  [`S0_NUMBER*AXI_AW    +: 1*AXI_AW ];
    assign s0_axi_arlen    = axi_arlen   [`S0_NUMBER*8         +: 1*8      ];
    assign s0_axi_arsize   = axi_arsize  [`S0_NUMBER*3         +: 1*3      ];
    assign s0_axi_arburst  = axi_arburst [`S0_NUMBER*2         +: 1*2      ];
    assign s0_axi_arlock   = axi_arlock  [`S0_NUMBER           +: 1        ];
    assign s0_axi_arcache  = axi_arcache [`S0_NUMBER*4         +: 1*4      ];
    assign s0_axi_arprot   = axi_arprot  [`S0_NUMBER*3         +: 1*3      ];
    assign s0_axi_arvalid  = axi_arvalid [`S0_NUMBER           +: 1        ];
    assign s0_axi_arready  = axi_arready [`S0_NUMBER           +: 1        ];
    assign s0_axi_rid      = axi_rid     [`S0_NUMBER*8         +: 1*8      ];
    assign s0_axi_rdata    = axi_rdata   [`S0_NUMBER*AXI_DW    +: 1*AXI_DW ];
    assign s0_axi_rresp    = axi_rresp   [`S0_NUMBER*2         +: 1*2      ];
    assign s0_axi_rlast    = axi_rlast   [`S0_NUMBER           +: 1        ];
    assign s0_axi_rvalid   = axi_rvalid  [`S0_NUMBER           +: 1        ];
    assign s0_axi_rready   = axi_rready  [`S0_NUMBER           +: 1        ];
    assign s1_axi_awid     = axi_awid    [`S1_NUMBER*8         +: 1*8      ];
    assign s1_axi_awaddr   = axi_awaddr  [`S1_NUMBER*AXI_AW    +: 1*AXI_AW ];
    assign s1_axi_awlen    = axi_awlen   [`S1_NUMBER*8         +: 1*8      ];
    assign s1_axi_awsize   = axi_awsize  [`S1_NUMBER*3         +: 1*3      ];
    assign s1_axi_awburst  = axi_awburst [`S1_NUMBER*2         +: 1*2      ];
    assign s1_axi_awlock   = axi_awlock  [`S1_NUMBER           +: 1        ];
    assign s1_axi_awcache  = axi_awcache [`S1_NUMBER*4         +: 1*4      ];
    assign s1_axi_awprot   = axi_awprot  [`S1_NUMBER*3         +: 1*3      ];
    assign s1_axi_awvalid  = axi_awvalid [`S1_NUMBER           +: 1        ];
    assign s1_axi_awready  = axi_awready [`S1_NUMBER           +: 1        ];
    assign s1_axi_wdata    = axi_wdata   [`S1_NUMBER*AXI_DW    +: 1*AXI_DW ];
    assign s1_axi_wstrb    = axi_wstrb   [`S1_NUMBER*AXI_SW    +: 1*AXI_SW ];
    assign s1_axi_wlast    = axi_wlast   [`S1_NUMBER           +: 1        ];
    assign s1_axi_wvalid   = axi_wvalid  [`S1_NUMBER           +: 1        ];
    assign s1_axi_wready   = axi_wready  [`S1_NUMBER           +: 1        ];
    assign s1_axi_bid      = axi_bid     [`S1_NUMBER*8         +: 1*8      ];
    assign s1_axi_bresp    = axi_bresp   [`S1_NUMBER*2         +: 1*2      ];
    assign s1_axi_bvalid   = axi_bvalid  [`S1_NUMBER           +: 1        ];
    assign s1_axi_bready   = axi_bready  [`S1_NUMBER           +: 1        ];
    assign s1_axi_arid     = axi_arid    [`S1_NUMBER*8         +: 1*8      ];
    assign s1_axi_araddr   = axi_araddr  [`S1_NUMBER*AXI_AW    +: 1*AXI_AW ];
    assign s1_axi_arlen    = axi_arlen   [`S1_NUMBER*8         +: 1*8      ];
    assign s1_axi_arsize   = axi_arsize  [`S1_NUMBER*3         +: 1*3      ];
    assign s1_axi_arburst  = axi_arburst [`S1_NUMBER*2         +: 1*2      ];
    assign s1_axi_arlock   = axi_arlock  [`S1_NUMBER           +: 1        ];
    assign s1_axi_arcache  = axi_arcache [`S1_NUMBER*4         +: 1*4      ];
    assign s1_axi_arprot   = axi_arprot  [`S1_NUMBER*3         +: 1*3      ];
    assign s1_axi_arvalid  = axi_arvalid [`S1_NUMBER           +: 1        ];
    assign s1_axi_arready  = axi_arready [`S1_NUMBER           +: 1        ];
    assign s1_axi_rid      = axi_rid     [`S1_NUMBER*8         +: 1*8      ];
    assign s1_axi_rdata    = axi_rdata   [`S1_NUMBER*AXI_DW    +: 1*AXI_DW ];
    assign s1_axi_rresp    = axi_rresp   [`S1_NUMBER*2         +: 1*2      ];
    assign s1_axi_rlast    = axi_rlast   [`S1_NUMBER           +: 1        ];
    assign s1_axi_rvalid   = axi_rvalid  [`S1_NUMBER           +: 1        ];
    assign s1_axi_rready   = axi_rready  [`S1_NUMBER           +: 1        ];    
    axi_ram #(
        .DATA_WIDTH                         (AXI_DW                    ),
        .ADDR_WIDTH                         (AXI_AW                    ),
        .ID_WIDTH                           (AXI_ID_WIDTH              ),
        .PIPELINE_OUTPUT                    (0                         ) 
    ) u_axi_ram (
        .clk                                (axi_aclk                 ),
        .rst                                (!axi_aresetn              ),
        .s_axi_awid                         (m0_axi_awid               ),
        .s_axi_awaddr                       (m0_axi_awaddr             ),
        .s_axi_awlen                        (m0_axi_awlen              ),
        .s_axi_awsize                       (m0_axi_awsize             ),
        .s_axi_awburst                      (m0_axi_awburst            ),
        .s_axi_awlock                       (m0_axi_awlock             ),
        .s_axi_awcache                      (m0_axi_awcache            ),
        .s_axi_awprot                       (m0_axi_awprot             ),
        .s_axi_awvalid                      (m0_axi_awvalid            ),
        .s_axi_awready                      (m0_axi_awready            ),
        .s_axi_wdata                        (m0_axi_wdata              ),
        .s_axi_wstrb                        (m0_axi_wstrb              ),
        .s_axi_wlast                        (m0_axi_wlast              ),
        .s_axi_wvalid                       (m0_axi_wvalid             ),
        .s_axi_wready                       (m0_axi_wready             ),
        .s_axi_bid                          (m0_axi_bid                ),
        .s_axi_bresp                        (m0_axi_bresp              ),
        .s_axi_bvalid                       (m0_axi_bvalid             ),
        .s_axi_bready                       (m0_axi_bready             ),
        .s_axi_arid                         (m0_axi_arid               ),
        .s_axi_araddr                       (m0_axi_araddr             ),
        .s_axi_arlen                        (m0_axi_arlen              ),
        .s_axi_arsize                       (m0_axi_arsize             ),
        .s_axi_arburst                      (m0_axi_arburst            ),
        .s_axi_arlock                       (m0_axi_arlock             ),
        .s_axi_arcache                      (m0_axi_arcache            ),
        .s_axi_arprot                       (m0_axi_arprot             ),
        .s_axi_arvalid                      (m0_axi_arvalid            ),
        .s_axi_arready                      (m0_axi_arready            ),
        .s_axi_rid                          (m0_axi_rid                ),
        .s_axi_rdata                        (m0_axi_rdata              ),
        .s_axi_rresp                        (m0_axi_rresp              ),
        .s_axi_rlast                        (m0_axi_rlast              ),
        .s_axi_rvalid                       (m0_axi_rvalid             ),
        .s_axi_rready                       (m0_axi_rready             ) 
    );
    axi_interconnect #(
        .S_COUNT   (S_COUNT),
        .M_COUNT   (M_COUNT),
        .DATA_WIDTH(AXI_DW),
        .ADDR_WIDTH(AXI_AW),
        .ID_WIDTH  (AXI_ID_WIDTH)
    ) u_axi_interconnect (
        .clk          (axi_aclk),
        .rst          (!axi_aresetn),
        //AXI slave interfaces
        .s_axi_awid   ({s1_axi_awid    , s0_axi_awid    }),
        .s_axi_awaddr ({s1_axi_awaddr  , s0_axi_awaddr  }),
        .s_axi_awlen  ({s1_axi_awlen   , s0_axi_awlen   }),
        .s_axi_awsize ({s1_axi_awsize  , s0_axi_awsize  }),
        .s_axi_awburst({s1_axi_awburst , s0_axi_awburst }),
        .s_axi_awlock ({s1_axi_awlock  , s0_axi_awlock  }),
        .s_axi_awcache({s1_axi_awcache , s0_axi_awcache }),
        .s_axi_awprot ({s1_axi_awprot  , s0_axi_awprot  }),
        .s_axi_awvalid({s1_axi_awvalid , s0_axi_awvalid }),
        .s_axi_awready({s1_axi_awready , s0_axi_awready }),
        .s_axi_wdata  ({s1_axi_wdata   , s0_axi_wdata   }),
        .s_axi_wstrb  ({s1_axi_wstrb   , s0_axi_wstrb   }),
        .s_axi_wlast  ({s1_axi_wlast   , s0_axi_wlast   }),
        .s_axi_wvalid ({s1_axi_wvalid  , s0_axi_wvalid  }),
        .s_axi_wready ({s1_axi_wready  , s0_axi_wready  }),
        .s_axi_bid    ({s1_axi_bid     , s0_axi_bid     }),
        .s_axi_bresp  ({s1_axi_bresp   , s0_axi_bresp   }),
        .s_axi_bvalid ({s1_axi_bvalid  , s0_axi_bvalid  }),
        .s_axi_bready ({s1_axi_bready  , s0_axi_bready  }),
        .s_axi_arid   ({s1_axi_arid    , s0_axi_arid    }),
        .s_axi_araddr ({s1_axi_araddr  , s0_axi_araddr  }),
        .s_axi_arlen  ({s1_axi_arlen   , s0_axi_arlen   }),
        .s_axi_arsize ({s1_axi_arsize  , s0_axi_arsize  }),
        .s_axi_arburst({s1_axi_arburst , s0_axi_arburst }),
        .s_axi_arlock ({s1_axi_arlock  , s0_axi_arlock  }),
        .s_axi_arcache({s1_axi_arcache , s0_axi_arcache }),
        .s_axi_arprot ({s1_axi_arprot  , s0_axi_arprot  }),
        .s_axi_arvalid({s1_axi_arvalid , s0_axi_arvalid }),
        .s_axi_arready({s1_axi_arready , s0_axi_arready }),
        .s_axi_rid    ({s1_axi_rid     , s0_axi_rid     }),
        .s_axi_rdata  ({s1_axi_rdata   , s0_axi_rdata   }),
        .s_axi_rresp  ({s1_axi_rresp   , s0_axi_rresp   }),
        .s_axi_rlast  ({s1_axi_rlast   , s0_axi_rlast   }),
        .s_axi_rvalid ({s1_axi_rvalid  , s0_axi_rvalid  }),
        .s_axi_rready ({s1_axi_rready  , s0_axi_rready  }),
        //AXI master interfaces
        .m_axi_awid   (m0_axi_awid                       ),//(axi_awid[2*8+:1*8]),
        .m_axi_awaddr (m0_axi_awaddr                     ),//(axi_awaddr[2*AXI_AW+:1*AXI_AW]),
        .m_axi_awlen  (m0_axi_awlen                      ),//(axi_awlen[2*8+:1*8]),
        .m_axi_awsize (m0_axi_awsize                     ),//(axi_awsize[2*3+:1*3]),
        .m_axi_awburst(m0_axi_awburst                    ),//(axi_awburst[2*2+:1*2]),
        .m_axi_awlock (m0_axi_awlock                     ),//(axi_awlock[2*1+:1*1]),
        .m_axi_awcache(m0_axi_awcache                    ),//(axi_awcache[2*4+:1*4]),
        .m_axi_awprot (m0_axi_awprot                     ),//(axi_awprot[2*3+:1*3]),
        .m_axi_awvalid(m0_axi_awvalid                    ),//(axi_awvalid[2*1+:1*1]),
        .m_axi_awready(m0_axi_awready                    ),//(axi_awready[2*1+:1*1]),
        .m_axi_wdata  (m0_axi_wdata                      ),//(axi_wdata[2*AXI_DW+:1*AXI_DW]),
        .m_axi_wstrb  (m0_axi_wstrb                      ),//(axi_wstrb[2*AXI_SW+:1*AXI_SW]),
        .m_axi_wlast  (m0_axi_wlast                      ),//(axi_wlast[2*1+:1*1]),
        .m_axi_wvalid (m0_axi_wvalid                     ),//(axi_wvalid[2*1+:1*1]),
        .m_axi_wready (m0_axi_wready                     ),//(axi_wready[2*1+:1*1]),
        .m_axi_bid    (m0_axi_bid                        ),//(axi_bid[2*8+:1*8]),
        .m_axi_bresp  (m0_axi_bresp                      ),//(axi_bresp[2*2+:1*2]),
        .m_axi_bvalid (m0_axi_bvalid                     ),//(axi_bvalid[2*1+:1*1]),
        .m_axi_bready (m0_axi_bready                     ),//(axi_bready[2*1+:1*1]),
        .m_axi_arid   (m0_axi_arid                       ),//(axi_arid[2*8+:1*8]),
        .m_axi_araddr (m0_axi_araddr                     ),//(axi_araddr[2*AXI_AW+:1*AXI_AW]),
        .m_axi_arlen  (m0_axi_arlen                      ),//(axi_arlen[2*8+:1*8]),
        .m_axi_arsize (m0_axi_arsize                     ),//(axi_arsize[2*3+:1*3]),
        .m_axi_arburst(m0_axi_arburst                    ),//(axi_arburst[2*2+:1*2]),
        .m_axi_arlock (m0_axi_arlock                     ),//(axi_arlock[2*1+:1*1]),
        .m_axi_arcache(m0_axi_arcache                    ),//(axi_arcache[2*4+:1*4]),
        .m_axi_arprot (m0_axi_arprot                     ),//(axi_arprot[2*3+:1*3]),
        .m_axi_arvalid(m0_axi_arvalid                    ),//(axi_arvalid[2*1+:1*1]),
        .m_axi_arready(m0_axi_arready                    ),//(axi_arready[2*1+:1*1]),
        .m_axi_rid    (m0_axi_rid                        ),//(axi_rid[2*8+:1*8]),
        .m_axi_rdata  (m0_axi_rdata                      ),//(axi_rdata[2*AXI_DW+:1*AXI_DW]),
        .m_axi_rresp  (m0_axi_rresp                      ),//(axi_rresp[2*2+:1*2]),
        .m_axi_rlast  (m0_axi_rlast                      ),//(axi_rlast[2*1+:1*1]),
        .m_axi_rvalid (m0_axi_rvalid                     ),//(axi_rvalid[2*1+:1*1]),
        .m_axi_rready (m0_axi_rready                     )//(axi_rready[2*1+:1*1])
    );
    //**********************************************************************************************
    image_to_ddr # (
        .CW                                 (CW                        ),
        .DW                                 (DW                        ),
        .AXI_AW                             (AXI_AW                    ),
        .IMAGE_WIDTH                        (IMAGE_WIDTH               ),
        .IMAGE_HEIGHT                       (IMAGE_HEIGHT              ) 
      )
      image0_to_ddr_inst (
        .i_Sys_clk                          (i_Sys_clk                 ),
        .i_Rst_n                            (i_Rst_n                   ),
        .i_Fix_en                           (1'b0                      ),
        .i_Din_field_sync                   (v_valid                   ),
        .i_Din_valid                        (h_valid                   ),
        .i_Din                              ({4'd0,hcnt}),//data_tmp                  ),
        .i_last_addr1                       ('d0                       ),
        .i_last_addr2                       ('d655360                  ),
        .o_last_wr_rst                      (user0_wr_rst              ),
        .o_last_wr_vs                       (user0_wr_vs               ),
        .o_last_wr_hs                       (user0_wr_hs               ),
        .o_last_wr_data                     (user0_wr_data             ),
        .o_last_wr_addr                     (user0_wr_axi_addr         ) 
      );    
      ddr_to_logic # (
        .CW                                 (CW                        ),
        .DW                                 (DW                        ),
        .AXI_AW                             (AXI_AW                    ),
        .IMAGE_WIDTH                        (IMAGE_WIDTH               ),
        .IMAGE_HEIGHT                       (IMAGE_HEIGHT              ) 
      )
      ddr_to_logic_inst (
        .i_Sys_clk                          (i_Sys_clk                 ),
        .i_Rst_n                            (i_Rst_n                   ),
        .i_Din_vs                           (v_valid               ),
        .i_Din_hs                           (h_valid               ),
        .i_last_addr1                       ('d0                       ),
        .i_last_addr2                       ('d655360                  ),
        .o_last_rd_rst                      (user0_rd_rst              ),
        .o_last_rd_vs                       (user0_rd_vs               ),
        .o_last_rd_hs                       (user0_rd_hs               ),
        .i_last_rd_data                     (user0_rd_data             ),
        .o_last_rd_addr                     (user0_rd_axi_addr         ),
        .o_Dout_valid                       (                          ),
        .o_Dout                             (                          ) 
      );      
    video_fdma # (
        .AXI_ID_DW                          (8                         ),
        .AXI_ID                             (0                         ),
        .AXI_AW                             (AXI_AW                    ),
        .AXI_DW                             (AXI_DW                    ),
        .DVP_DATA_WIDTH                     (DVP_DATA_WIDTH            ) 
      )
      video0_fdma_inst (
        .dvp_wr_rst                         (user0_wr_rst                ),
        .dvp_wr_clk                         (user0_wr_clk                ),
        .dvp_wr_vs                          (user0_wr_vs                 ),
        .dvp_wr_hs                          (user0_wr_hs                 ),
        .dvp_wr_data                        (user0_wr_data               ),
        .dvp_wr_axi_addr                    (user0_wr_axi_addr           ),

        .dvp_rd_rst                         (user0_rd_rst                ),
        .dvp_rd_clk                         (user0_rd_clk                ),
        .dvp_rd_vs                          (user0_rd_vs                 ),
        .dvp_rd_hs                          (user0_rd_hs                 ),
        .dvp_rd_data_valid                  (user0_rd_data_valid         ),
        .dvp_rd_data                        (user0_rd_data               ),
        .dvp_rd_axi_addr                    (user0_rd_axi_addr           ),
        .clk_axi                         (axi_aclk                   ),
        .rst_axi                      (~axi_aresetn                ),
        .m_axi_awid                         (s0_axi_awid                ),
        .m_axi_awaddr                       (s0_axi_awaddr              ),
        .m_axi_awlen                        (s0_axi_awlen               ),
        .m_axi_awsize                       (s0_axi_awsize              ),
        .m_axi_awburst                      (s0_axi_awburst             ),
        .m_axi_awlock                       (s0_axi_awlock              ),
        .m_axi_awcache                      (s0_axi_awcache             ),
        .m_axi_awprot                       (s0_axi_awprot              ),
        // .m_axi_awqos                        (s0_axi_awqos               ),
        .m_axi_awvalid                      (s0_axi_awvalid             ),
        .m_axi_awready                      (s0_axi_awready             ),
        // .m_axi_wid                          (s0_axi_wid                 ),
        .m_axi_wdata                        (s0_axi_wdata               ),
        .m_axi_wstrb                        (s0_axi_wstrb               ),
        .m_axi_wlast                        (s0_axi_wlast               ),
        .m_axi_wvalid                       (s0_axi_wvalid              ),
        .m_axi_wready                       (s0_axi_wready              ),
        .m_axi_bid                          (s0_axi_bid                 ),
        .m_axi_bresp                        (s0_axi_bresp               ),
        .m_axi_bvalid                       (s0_axi_bvalid              ),
        .m_axi_bready                       (s0_axi_bready              ),
        .m_axi_arid                         (s0_axi_arid                ),
        .m_axi_araddr                       (s0_axi_araddr              ),
        .m_axi_arlen                        (s0_axi_arlen               ),
        .m_axi_arsize                       (s0_axi_arsize              ),
        .m_axi_arburst                      (s0_axi_arburst             ),
        .m_axi_arlock                       (s0_axi_arlock              ),
        .m_axi_arcache                      (s0_axi_arcache             ),
        .m_axi_arprot                       (s0_axi_arprot              ),
        // .m_axi_arqos                        (s0_axi_arqos               ),
        .m_axi_arvalid                      (s0_axi_arvalid             ),
        .m_axi_arready                      (s0_axi_arready             ),
        .m_axi_rid                          (s0_axi_rid                 ),
        .m_axi_rdata                        (s0_axi_rdata               ),
        .m_axi_rresp                        (s0_axi_rresp               ),
        .m_axi_rlast                        (s0_axi_rlast               ),
        .m_axi_rvalid                       (s0_axi_rvalid              ),
        .m_axi_rready                       (s0_axi_rready              ) 
      );    
    //**********************************************************************************************
    // image_to_ddr # (
    //     .CW                                 (CW                        ),
    //     .DW                                 (DW                        ),
    //     .AXI_AW                             (AXI_AW                    ),
    //     .IMAGE_WIDTH                        (IMAGE_WIDTH               ),
    //     .IMAGE_HEIGHT                       (IMAGE_HEIGHT              ) 
    //   )
    //   image1_to_ddr_inst (
    //     .i_Sys_clk                          (i_Sys_clk                 ),
    //     .i_Rst_n                            (i_Rst_n                   ),
    //     .i_Fix_en                           (1'b0                      ),
    //     .i_Din_field_sync                        (v_valid                   ),
    //     .i_Din_valid                        (h_valid                   ),
    //     .i_Din                              ({4'd0,hcnt}),//data_tmp                  ),
    //     .i_last_addr1                       ('d0                       ),
    //     .i_last_addr2                       ('d0                       ),
    //     .o_last_wr_rst                      (user1_wr_rst              ),
    //     .o_last_wr_vs                      (user1_wr_vs              ),
    //     .o_last_wr_hs                      (user1_wr_hs               ),
    //     .o_last_wr_data                     (user1_wr_data             ),
    //     .o_last_wr_addr                     (user1_wr_axi_addr         ) 
    //   );    
    //   video_fdma # (
    //     .AXI_ID_DW                          (8                         ),
    //     .AXI_ID                             (1                         ),
    //     .AXI_AW                             (AXI_AW                    ),
    //     .AXI_DW                             (AXI_DW                    ),
    //     .DVP_DATA_WIDTH                     (DVP_DATA_WIDTH            ) 
    //   )
    //   video1_fdma_inst (
    //     .dvp_wr_rst                         (user1_wr_rst                ),
    //     .dvp_wr_clk                         (user1_wr_clk                ),
    //     .dvp_wr_vs                          (user1_wr_vs                 ),
    //     .dvp_wr_hs                          (user1_wr_hs                 ),
    //     .dvp_wr_data                        (user1_wr_data               ),
    //     .dvp_wr_axi_addr                    (user1_wr_axi_addr           ),
    //     .dvp_rd_rst                         (user1_rd_rst                ),
    //     .dvp_rd_clk                         (user1_rd_clk                ),
    //     .dvp_rd_vs                          (user1_rd_vs                 ),
    //     .dvp_rd_hs                          (user1_rd_hs                 ),
    //     .dvp_rd_data_valid                  (user1_rd_data_valid         ),
    //     .dvp_rd_data                        (user1_rd_data               ),
    //     .dvp_rd_axi_addr                    (user1_rd_axi_addr           ),
    //     .clk_axi                         (axi_aclk                ),
    //     .rst_axi                      (~axi_aresetn             ),
    //     .m_axi_awid                         (s1_axi_awid                ),
    //     .m_axi_awaddr                       (s1_axi_awaddr              ),
    //     .m_axi_awlen                        (s1_axi_awlen               ),
    //     .m_axi_awsize                       (s1_axi_awsize              ),
    //     .m_axi_awburst                      (s1_axi_awburst             ),
    //     .m_axi_awlock                       (s1_axi_awlock              ),
    //     .m_axi_awcache                      (s1_axi_awcache             ),
    //     .m_axi_awprot                       (s1_axi_awprot              ),
    //     // .m_axi_awqos                        (s1_axi_awqos               ),
    //     .m_axi_awvalid                      (s1_axi_awvalid             ),
    //     .m_axi_awready                      (s1_axi_awready             ),
    //     // .m_axi_wid                          (s1_axi_wid                 ),
    //     .m_axi_wdata                        (s1_axi_wdata               ),
    //     .m_axi_wstrb                        (s1_axi_wstrb               ),
    //     .m_axi_wlast                        (s1_axi_wlast               ),
    //     .m_axi_wvalid                       (s1_axi_wvalid              ),
    //     .m_axi_wready                       (s1_axi_wready              ),
    //     .m_axi_bid                          (s1_axi_bid                 ),
    //     .m_axi_bresp                        (s1_axi_bresp               ),
    //     .m_axi_bvalid                       (s1_axi_bvalid              ),
    //     .m_axi_bready                       (s1_axi_bready              ),
    //     .m_axi_arid                         (s1_axi_arid                ),
    //     .m_axi_araddr                       (s1_axi_araddr              ),
    //     .m_axi_arlen                        (s1_axi_arlen               ),
    //     .m_axi_arsize                       (s1_axi_arsize              ),
    //     .m_axi_arburst                      (s1_axi_arburst             ),
    //     .m_axi_arlock                       (s1_axi_arlock              ),
    //     .m_axi_arcache                      (s1_axi_arcache             ),
    //     .m_axi_arprot                       (s1_axi_arprot              ),
    //     // .m_axi_arqos                        (s1_axi_arqos               ),
    //     .m_axi_arvalid                      (s1_axi_arvalid             ),
    //     .m_axi_arready                      (s1_axi_arready             ),
    //     .m_axi_rid                          (s1_axi_rid                 ),
    //     .m_axi_rdata                        (s1_axi_rdata               ),
    //     .m_axi_rresp                        (s1_axi_rresp               ),
    //     .m_axi_rlast                        (s1_axi_rlast               ),
    //     .m_axi_rvalid                       (s1_axi_rvalid              ),
    //     .m_axi_rready                       (s1_axi_rready              ) 
    //   );      
    //**********************************************************************************************
endmodule

