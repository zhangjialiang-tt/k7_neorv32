-- megafunction wizard: %RAM: 2-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram

-- ============================================================
-- File Name: lpm_dual_clk_port_ram.vhd
-- Megafunction Name(s):
-- 			altsyncram
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 17.0.0 Build 595 04/25/2017 SJ Standard Edition
-- ************************************************************


--Copyright (C) 2017  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions
--and other software and tools, and its AMPP partner logic
--functions, and any output files from any of the foregoing
--(including device programming or simulation files), and any
--associated documentation or information are expressly subject
--to the terms and conditions of the Intel Program License
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel MegaCore Function License Agreement, or other
--applicable license agreement, including, without limitation,
--that your use is for the sole purpose of programming logic
--devices manufactured by Intel and sold by Intel or its
--authorized distributors.  Please refer to the applicable
--agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

-- LIBRARY altera_mf;
-- USE altera_mf.altera_mf_components.all;

ENTITY lpm_dual_clk_port_ram IS
    generic
    (
        DATA_WIDTH        : integer := 16;            --data width
        ADDR_WIDTH        : integer := 10;            --addr width
        ADDR_DEPTH        : integer := 1024           --
    );
    PORT
    (
        address_a     : IN STD_LOGIC_VECTOR (ADDR_WIDTH - 1 DOWNTO 0);
        address_b     : IN STD_LOGIC_VECTOR (ADDR_WIDTH - 1 DOWNTO 0);
        clock_a       : IN STD_LOGIC  := '1';
        clock_b       : IN STD_LOGIC ;
        data_a        : IN STD_LOGIC_VECTOR (DATA_WIDTH - 1 DOWNTO 0);
        data_b        : IN STD_LOGIC_VECTOR (DATA_WIDTH - 1 DOWNTO 0);
        enable_a      : IN STD_LOGIC  := '1';
        enable_b      : IN STD_LOGIC  := '1';
        rden_a        : IN STD_LOGIC  := '1';
        rden_b        : IN STD_LOGIC  := '1';
        wren_a        : IN STD_LOGIC  := '0';
        wren_b        : IN STD_LOGIC  := '0';
        q_a           : OUT STD_LOGIC_VECTOR (DATA_WIDTH - 1 DOWNTO 0);
        q_b           : OUT STD_LOGIC_VECTOR (DATA_WIDTH - 1 DOWNTO 0)
    );
END lpm_dual_clk_port_ram;


ARCHITECTURE SYN OF lpm_dual_clk_port_ram IS

COMPONENT true_dual_port_ram
generic
(
DATA_WIDTH      : NATURAL  := 8;
ADDR_WIDTH      : NATURAL  := 9;
WRITE_MODE_1    : STRING   := "READ_FIRST";	-- WRITE_FIRST; READ_FIRST; NO_CHANGE
WRITE_MODE_2    : STRING   := "READ_FIRST";
OUTPUT_REG_1    : STRING   := "FALSE";
OUTPUT_REG_2    : STRING   := "FALSE";
RAM_INIT_FILE   : STRING   := "ram_init_file.mem"
);
PORT
(
we1             :  in  std_logic  ;
we2             :  in  std_logic  ;
clka            :  in  std_logic  ;
clkb            :  in  std_logic  ;
din1            :  in  std_logic_vector(DATA_WIDTH-1 downto 0)  ;
din2            :  in  std_logic_vector(DATA_WIDTH-1 downto 0)  ;
addr1           :  in  std_logic_vector(ADDR_WIDTH-1 downto 0)  ;
addr2           :  in  std_logic_vector(ADDR_WIDTH-1 downto 0)  ;
dout1           :  out std_logic_vector(DATA_WIDTH-1 downto 0)  ;
dout2           :  out std_logic_vector(DATA_WIDTH-1 downto 0)
);
END COMPONENT;

    signal write_enable_1 : std_logic;
    signal write_enable_2 : std_logic;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (DATA_WIDTH - 1 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (DATA_WIDTH - 1 DOWNTO 0);

BEGIN
	q_a    <= sub_wire0(DATA_WIDTH - 1 DOWNTO 0);
	q_b    <= sub_wire1(DATA_WIDTH - 1 DOWNTO 0);

--  	altsyncram_component : altsyncram
--  	GENERIC MAP
--  	(
--  		address_reg_b => "CLOCK1",
--  		clock_enable_input_a => "NORMAL",
--  		clock_enable_input_b => "NORMAL",
--  		clock_enable_output_a => "BYPASS",
--  		clock_enable_output_b => "BYPASS",
--  		indata_reg_b => "CLOCK1",
--  		intended_device_family => "CYCLONE IV E",
--  		lpm_type => "altsyncram",
--  		numwords_a => ADDR_DEPTH,
--  		numwords_b => ADDR_DEPTH,
--  		operation_mode => "BIDIR_DUAL_PORT",
--  		outdata_aclr_a => "NONE",
--  		outdata_aclr_b => "NONE",
--  		outdata_reg_a => "UNREGISTERED",
--  		outdata_reg_b => "UNREGISTERED",
--  		power_up_uninitialized => "FALSE",
--  		read_during_write_mode_mixed_ports => "DONT_CARE",
--  		read_during_write_mode_port_a => "NEW_DATA_NO_NBE_READ",
--  		read_during_write_mode_port_b => "NEW_DATA_NO_NBE_READ",
--  		widthad_a => ADDR_WIDTH,
--  		widthad_b => ADDR_WIDTH,
--  		width_a => DATA_WIDTH,
--  		width_b => DATA_WIDTH,
--  		width_byteena_a => 1,
--  		width_byteena_b => 1,
--  		wrcontrol_wraddress_reg_b => "CLOCK1"
--  	)
--  	PORT MAP
--  	(
--  		address_a => address_a,
--  		address_b => address_b,
--  		clock0    => clock_a,
--  		clock1    => clock_b,
--  		clocken0  => enable_a,
--  		clocken1  => enable_b,
--  		data_a    => data_a,
--  		data_b    => data_b,
--  		rden_a    => rden_a,
--  		rden_b    => rden_b,
--  		wren_a    => wren_a,
--  		wren_b    => wren_b,
--  		q_a       => sub_wire0,
--  		q_b       => sub_wire1
--  	);

    write_enable_1 <= (enable_a and wren_a);
    write_enable_2 <= (enable_b and wren_b);

    altsyncram_component : true_dual_port_ram
    generic map
    (
        DATA_WIDTH      => DATA_WIDTH,
        ADDR_WIDTH      => ADDR_WIDTH,
        WRITE_MODE_1    => "READ_FIRST",
        WRITE_MODE_2    => "READ_FIRST",
        OUTPUT_REG_1    => "FALSE",
        OUTPUT_REG_2    => "FALSE",
        RAM_INIT_FILE   => "ram_init_file.mem"
    )
    PORT map
    (
        we1             => write_enable_1,
        we2             => write_enable_2,
        clka            => clock_a,
        clkb            => clock_b,
        din1            => data_a,
        din2            => data_b,
        addr1           => address_a,
        addr2           => address_b,
        dout1           => sub_wire0,
        dout2           => sub_wire1
    );


END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ADDRESSSTALL_A NUMERIC "0"
-- Retrieval info: PRIVATE: ADDRESSSTALL_B NUMERIC "0"
-- Retrieval info: PRIVATE: BYTEENA_ACLR_A NUMERIC "0"
-- Retrieval info: PRIVATE: BYTEENA_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_ENABLE_A NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_ENABLE_B NUMERIC "0"
-- Retrieval info: PRIVATE: BYTE_SIZE NUMERIC "8"
-- Retrieval info: PRIVATE: BlankMemory NUMERIC "1"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_A NUMERIC "1"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_INPUT_B NUMERIC "1"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_OUTPUT_A NUMERIC "1"
-- Retrieval info: PRIVATE: CLOCK_ENABLE_OUTPUT_B NUMERIC "1"
-- Retrieval info: PRIVATE: CLRdata NUMERIC "0"
-- Retrieval info: PRIVATE: CLRq NUMERIC "0"
-- Retrieval info: PRIVATE: CLRrdaddress NUMERIC "0"
-- Retrieval info: PRIVATE: CLRrren NUMERIC "0"
-- Retrieval info: PRIVATE: CLRwraddress NUMERIC "0"
-- Retrieval info: PRIVATE: CLRwren NUMERIC "0"
-- Retrieval info: PRIVATE: Clock NUMERIC "5"
-- Retrieval info: PRIVATE: Clock_A NUMERIC "0"
-- Retrieval info: PRIVATE: Clock_B NUMERIC "0"
-- Retrieval info: PRIVATE: IMPLEMENT_IN_LES NUMERIC "0"
-- Retrieval info: PRIVATE: INDATA_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: INDATA_REG_B NUMERIC "1"
-- Retrieval info: PRIVATE: INIT_FILE_LAYOUT STRING "PORT_A"
-- Retrieval info: PRIVATE: INIT_TO_SIM_X NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "MAX 10"
-- Retrieval info: PRIVATE: JTAG_ENABLED NUMERIC "0"
-- Retrieval info: PRIVATE: JTAG_ID STRING "NONE"
-- Retrieval info: PRIVATE: MAXIMUM_DEPTH NUMERIC "0"
-- Retrieval info: PRIVATE: MEMSIZE NUMERIC "16384"
-- Retrieval info: PRIVATE: MEM_IN_BITS NUMERIC "0"
-- Retrieval info: PRIVATE: MIFfilename STRING ""
-- Retrieval info: PRIVATE: OPERATION_MODE NUMERIC "3"
-- Retrieval info: PRIVATE: OUTDATA_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: OUTDATA_REG_B NUMERIC "0"
-- Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
-- Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_MIXED_PORTS NUMERIC "2"
-- Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_PORT_A NUMERIC "4"
-- Retrieval info: PRIVATE: READ_DURING_WRITE_MODE_PORT_B NUMERIC "4"
-- Retrieval info: PRIVATE: REGdata NUMERIC "1"
-- Retrieval info: PRIVATE: REGq NUMERIC "0"
-- Retrieval info: PRIVATE: REGrdaddress NUMERIC "0"
-- Retrieval info: PRIVATE: REGrren NUMERIC "1"
-- Retrieval info: PRIVATE: REGwraddress NUMERIC "1"
-- Retrieval info: PRIVATE: REGwren NUMERIC "1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: USE_DIFF_CLKEN NUMERIC "0"
-- Retrieval info: PRIVATE: UseDPRAM NUMERIC "1"
-- Retrieval info: PRIVATE: VarWidth NUMERIC "0"
-- Retrieval info: PRIVATE: WIDTH_READ_A NUMERIC "16"
-- Retrieval info: PRIVATE: WIDTH_READ_B NUMERIC "16"
-- Retrieval info: PRIVATE: WIDTH_WRITE_A NUMERIC "16"
-- Retrieval info: PRIVATE: WIDTH_WRITE_B NUMERIC "16"
-- Retrieval info: PRIVATE: WRADDR_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: WRADDR_REG_B NUMERIC "1"
-- Retrieval info: PRIVATE: WRCTRL_ACLR_B NUMERIC "0"
-- Retrieval info: PRIVATE: enable NUMERIC "1"
-- Retrieval info: PRIVATE: rden NUMERIC "1"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: ADDRESS_REG_B STRING "CLOCK1"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_A STRING "NORMAL"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_INPUT_B STRING "NORMAL"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_OUTPUT_A STRING "BYPASS"
-- Retrieval info: CONSTANT: CLOCK_ENABLE_OUTPUT_B STRING "BYPASS"
-- Retrieval info: CONSTANT: INDATA_REG_B STRING "CLOCK1"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "MAX 10"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altsyncram"
-- Retrieval info: CONSTANT: NUMWORDS_A NUMERIC "1024"
-- Retrieval info: CONSTANT: NUMWORDS_B NUMERIC "1024"
-- Retrieval info: CONSTANT: OPERATION_MODE STRING "BIDIR_DUAL_PORT"
-- Retrieval info: CONSTANT: OUTDATA_ACLR_A STRING "NONE"
-- Retrieval info: CONSTANT: OUTDATA_ACLR_B STRING "NONE"
-- Retrieval info: CONSTANT: OUTDATA_REG_A STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: OUTDATA_REG_B STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: POWER_UP_UNINITIALIZED STRING "FALSE"
-- Retrieval info: CONSTANT: READ_DURING_WRITE_MODE_PORT_A STRING "NEW_DATA_WITH_NBE_READ"
-- Retrieval info: CONSTANT: READ_DURING_WRITE_MODE_PORT_B STRING "NEW_DATA_WITH_NBE_READ"
-- Retrieval info: CONSTANT: WIDTHAD_A NUMERIC "10"
-- Retrieval info: CONSTANT: WIDTHAD_B NUMERIC "10"
-- Retrieval info: CONSTANT: WIDTH_A NUMERIC "16"
-- Retrieval info: CONSTANT: WIDTH_B NUMERIC "16"
-- Retrieval info: CONSTANT: WIDTH_BYTEENA_A NUMERIC "1"
-- Retrieval info: CONSTANT: WIDTH_BYTEENA_B NUMERIC "1"
-- Retrieval info: CONSTANT: WRCONTROL_WRADDRESS_REG_B STRING "CLOCK1"
-- Retrieval info: USED_PORT: address_a 0 0 10 0 INPUT NODEFVAL "address_a[9..0]"
-- Retrieval info: USED_PORT: address_b 0 0 10 0 INPUT NODEFVAL "address_b[9..0]"
-- Retrieval info: USED_PORT: clock_a 0 0 0 0 INPUT VCC "clock_a"
-- Retrieval info: USED_PORT: clock_b 0 0 0 0 INPUT NODEFVAL "clock_b"
-- Retrieval info: USED_PORT: data_a 0 0 16 0 INPUT NODEFVAL "data_a[15..0]"
-- Retrieval info: USED_PORT: data_b 0 0 16 0 INPUT NODEFVAL "data_b[15..0]"
-- Retrieval info: USED_PORT: enable_a 0 0 0 0 INPUT VCC "enable_a"
-- Retrieval info: USED_PORT: enable_b 0 0 0 0 INPUT VCC "enable_b"
-- Retrieval info: USED_PORT: q_a 0 0 16 0 OUTPUT NODEFVAL "q_a[15..0]"
-- Retrieval info: USED_PORT: q_b 0 0 16 0 OUTPUT NODEFVAL "q_b[15..0]"
-- Retrieval info: USED_PORT: rden_a 0 0 0 0 INPUT VCC "rden_a"
-- Retrieval info: USED_PORT: rden_b 0 0 0 0 INPUT VCC "rden_b"
-- Retrieval info: USED_PORT: wren_a 0 0 0 0 INPUT GND "wren_a"
-- Retrieval info: USED_PORT: wren_b 0 0 0 0 INPUT GND "wren_b"
-- Retrieval info: CONNECT: @address_a 0 0 10 0 address_a 0 0 10 0
-- Retrieval info: CONNECT: @address_b 0 0 10 0 address_b 0 0 10 0
-- Retrieval info: CONNECT: @clock0 0 0 0 0 clock_a 0 0 0 0
-- Retrieval info: CONNECT: @clock1 0 0 0 0 clock_b 0 0 0 0
-- Retrieval info: CONNECT: @clocken0 0 0 0 0 enable_a 0 0 0 0
-- Retrieval info: CONNECT: @clocken1 0 0 0 0 enable_b 0 0 0 0
-- Retrieval info: CONNECT: @data_a 0 0 16 0 data_a 0 0 16 0
-- Retrieval info: CONNECT: @data_b 0 0 16 0 data_b 0 0 16 0
-- Retrieval info: CONNECT: @rden_a 0 0 0 0 rden_a 0 0 0 0
-- Retrieval info: CONNECT: @rden_b 0 0 0 0 rden_b 0 0 0 0
-- Retrieval info: CONNECT: @wren_a 0 0 0 0 wren_a 0 0 0 0
-- Retrieval info: CONNECT: @wren_b 0 0 0 0 wren_b 0 0 0 0
-- Retrieval info: CONNECT: q_a 0 0 16 0 @q_a 0 0 16 0
-- Retrieval info: CONNECT: q_b 0 0 16 0 @q_b 0 0 16 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_dual_clk_port_ram.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_dual_clk_port_ram.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_dual_clk_port_ram.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_dual_clk_port_ram.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_dual_clk_port_ram_inst.vhd TRUE
-- Retrieval info: LIB_FILE: altera_mf
