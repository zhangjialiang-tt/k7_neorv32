-- megafunction wizard: %lpm_mult%
-- generation: standard
-- version: wm1.0
-- module: lpm_mult

-- ============================================================
-- file name: multi_un_16x16.vhd
-- megafunction name(s):
-- 			lpm_mult
--
-- simulation library files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- this is a wizard-generated file. do not edit this file!
--
-- 13.1.4 build 182 03/12/2014 sj full version
-- ************************************************************


--copyright (c) 1991-2014 altera corporation
--your use of altera corporation's design tools, logic functions
--and other software and tools, and its ampp partner logic
--functions, and any output files from any of the foregoing
--(including device programming or simulation files), and any
--associated documentation or information are expressly subject
--to the terms and conditions of the altera program license
--subscription agreement, altera megacore function license
--agreement, or other applicable license agreement, including,
--without limitation, that your use is for the sole purpose of
--programming logic devices manufactured by altera and sold by
--altera or its authorized distributors.  please refer to the
--applicable agreement for further details.


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

--library lpm;
--use lpm.all;

entity multi_mxn is
    generic
    (
        LPM_PIPELINE        : natural;
        LPM_WIDTHA          : natural;
        LPM_WIDTHB          : natural;
        LPM_REPRESENTATION  : string;
        LPM_RESET_ENABLE	: NATURAL:=0
    );
    port
    (
        rst_n       : in std_logic :='0';
        clken		: in std_logic ;
        clock		: in std_logic ;
        dataa		: in std_logic_vector (LPM_WIDTHA - 1 downto 0);
        datab		: in std_logic_vector (LPM_WIDTHB - 1 downto 0);
        result		: out std_logic_vector (LPM_WIDTHA + LPM_WIDTHB - 1 downto 0)
    );
end multi_mxn;


architecture syn of multi_mxn is

signal dataa_tmp    : std_logic_vector   (LPM_WIDTHA-1 downto 0) ;
signal datab_tmp    : std_logic_vector   (LPM_WIDTHB-1 downto 0) ;
signal sub_wire0	: std_logic_vector (LPM_WIDTHA + LPM_WIDTHB - 1 downto 0);

signal reset_cnt    : unsigned (7 downto 0) := to_unsigned(0,8);
signal reset_n_inter: std_logic;
--  component lpm_mult
--  generic (
--      lpm_hint		: string;
--  		lpm_pipeline		: natural;
--  		lpm_representation		: string;
--  		lpm_type		: string;
--  		lpm_widtha		: natural;
--  		lpm_widthb		: natural;
--  		lpm_widthp		: natural
--      );
--  port (
--      aclr	: in std_logic ;
--      clock	: in std_logic ;
--      sum     : in std_logic;
--      datab	: in std_logic_vector (lpm_widthb - 1 downto 0);
--      clken	: in std_logic ;
--      dataa	: in std_logic_vector (lpm_widtha - 1 downto 0);
--      result	: out std_logic_vector (lpm_widthp - 1 downto 0)
--      );
--  end component;


component parallel_ppl_mult
generic
(
MUL1_WIDTH : natural := 36                      ;
MUL2_WIDTH : natural := 26                      ;
PPL_LEVEL  : natural := 5                       ;
SINED      : string  := "YES"                   ;
MUL_IREG   : string  := "YES"                   ;
PROD_WIDTH : natural := 62
);
port
(
clk        : in  std_logic                                  ;
rst_n      : in  std_logic                                  ;
mul1       : in  std_logic_vector   (MUL1_WIDTH-1 downto 0) ;
mul2       : in  std_logic_vector   (MUL2_WIDTH-1 downto 0) ;
prod       : out std_logic_vector   (PROD_WIDTH-1 downto 0)
);
end component;

begin

    result    <= sub_wire0(LPM_WIDTHA + LPM_WIDTHB - 1 downto 0);

--      lpm_mult_component : lpm_mult
--      generic map
--      (
--          lpm_hint            => "maximize_speed=5",
--        		lpm_pipeline        => LPM_PIPELINE,
--        		lpm_representation  => LPM_REPRESENTATION,
--        		lpm_type            => "lpm_mult",
--        		lpm_widtha          => LPM_WIDTHA,
--        		lpm_widthb          => LPM_WIDTHB,
--        		lpm_widthp          => LPM_WIDTHA + LPM_WIDTHB
--      )
--      port map
--      (
--          aclr => '0',
--          clock => clock,
--          datab => datab,
--          clken => clken,
--          dataa => dataa,
--          sum => '0',
--          result => sub_wire0
--      );

    LPM_RESET_ENABLE0 : if(LPM_RESET_ENABLE = 0)generate
        reset_n_inter   <=  '1' when (reset_cnt >= 198) else
                            '0';

        dataa_tmp       <=  dataa when (reset_cnt >= 100) else
                            (others => '0');
        datab_tmp       <=  datab when (reset_cnt >= 100) else
                            (others => '0');
    end generate;

    LPM_RESET_ENABLE1 : if(LPM_RESET_ENABLE = 1)generate
        reset_n_inter   <=  rst_n;
        dataa_tmp       <=  dataa ;
        datab_tmp       <=  datab ;
    end generate;


    process(clock)
    begin
        if(rising_edge(clock))then
            if (reset_cnt <  200) then
                reset_cnt <= reset_cnt + 1;
            end if;
        end if;
    end process;

    lpm_mult_component : parallel_ppl_mult
    generic map
    (
        PPL_LEVEL   => LPM_PIPELINE,
        SINED       => LPM_REPRESENTATION,
        MUL_IREG    => "YES",
        MUL1_WIDTH  => LPM_WIDTHA,
        MUL2_WIDTH  => LPM_WIDTHB,
        PROD_WIDTH  => LPM_WIDTHA + LPM_WIDTHB
    )
    port map
    (
        clk         => clock,
        rst_n       => reset_n_inter ,
        mul1        => dataa_tmp,
        mul2        => datab_tmp,
        prod        => sub_wire0
    );

end syn;
